module d1_mul_acc (
    input dense_sum_i,
    input dense_w_i,
    input dense_b_i,
    input dense_input_i,
    output dense_output_o
);



endmodule