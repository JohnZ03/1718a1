module dense_1 (
    clk,
    rst_n,
    
);
    
endmodule